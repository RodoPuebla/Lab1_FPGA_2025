LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Multiplicador_SS IS 
	PORT
	(
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		S0 :  OUT  STD_LOGIC;
		S1 :  OUT  STD_LOGIC;
		S2 :  OUT  STD_LOGIC;
		C1 :  OUT  STD_LOGIC
	);
END Multiplicador_SS;

ARCHITECTURE bdf_type OF Multiplicador_SS IS 

COMPONENT full_adder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 C_in : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 C_out : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_2 <= '0';
SYNTHESIZED_WIRE_4 <= '0';



S0 <= A0 AND B0;


b2v_inst2 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_0,
		 B => SYNTHESIZED_WIRE_1,
		 C_in => SYNTHESIZED_WIRE_2,
		 S => S1,
		 C_out => SYNTHESIZED_WIRE_5);


SYNTHESIZED_WIRE_1 <= B0 AND A1;



b2v_inst5 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_3,
		 B => SYNTHESIZED_WIRE_4,
		 C_in => SYNTHESIZED_WIRE_5,
		 S => S2,
		 C_out => C1);


SYNTHESIZED_WIRE_3 <= B1 AND A1;


SYNTHESIZED_WIRE_0 <= A0 AND B1;



END bdf_type;