LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Multiplicador_CS IS 
	PORT
	(
		A0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		S0 :  OUT  STD_LOGIC;
		S1 :  OUT  STD_LOGIC;
		S2 :  OUT  STD_LOGIC;
		C1 :  OUT  STD_LOGIC;
		Bandera_Z :  OUT  STD_LOGIC
	);
END Multiplicador_CS;

ARCHITECTURE bdf_type OF Multiplicador_CS IS 

COMPONENT full_adder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 C_in : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 C_out : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_37 <= '0';
SYNTHESIZED_WIRE_26 <= '0';
SYNTHESIZED_WIRE_28 <= '1';



SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_43 <= SYNTHESIZED_WIRE_35 AND SYNTHESIZED_WIRE_33;


b2v_inst10 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_36,
		 B => SYNTHESIZED_WIRE_37,
		 C_in => SYNTHESIZED_WIRE_2,
		 S => SYNTHESIZED_WIRE_3,
		 C_out => SYNTHESIZED_WIRE_6);


SYNTHESIZED_WIRE_39 <= SYNTHESIZED_WIRE_34 AND SYNTHESIZED_WIRE_33;


SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_3;


SYNTHESIZED_WIRE_36 <= NOT(SYNTHESIZED_WIRE_34);



b2v_inst14 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_36,
		 B => SYNTHESIZED_WIRE_37,
		 C_in => SYNTHESIZED_WIRE_6,
		 S => SYNTHESIZED_WIRE_10);


b2v_inst15 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_39,
		 B => SYNTHESIZED_WIRE_8,
		 C_in => SYNTHESIZED_WIRE_9,
		 S => SYNTHESIZED_WIRE_40);


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_10;


Bandera_Z <= SYNTHESIZED_WIRE_11 AND SYNTHESIZED_WIRE_12 AND SYNTHESIZED_WIRE_13 AND SYNTHESIZED_WIRE_14;


SYNTHESIZED_WIRE_11 <= NOT(SYNTHESIZED_WIRE_40);



SYNTHESIZED_WIRE_12 <= NOT(SYNTHESIZED_WIRE_41);




SYNTHESIZED_WIRE_13 <= NOT(SYNTHESIZED_WIRE_42);



SYNTHESIZED_WIRE_14 <= NOT(SYNTHESIZED_WIRE_43);



PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_35 <= A0;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_33 <= B0;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_38 <= B1;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_34 <= A1;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	S0 <= SYNTHESIZED_WIRE_43;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	S1 <= SYNTHESIZED_WIRE_42;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	C1 <= SYNTHESIZED_WIRE_40;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	S2 <= SYNTHESIZED_WIRE_41;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_23;



b2v_inst5 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_24,
		 B => SYNTHESIZED_WIRE_25,
		 C_in => SYNTHESIZED_WIRE_26,
		 S => SYNTHESIZED_WIRE_42,
		 C_out => SYNTHESIZED_WIRE_32);


b2v_inst6 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_27,
		 B => SYNTHESIZED_WIRE_28,
		 C_in => SYNTHESIZED_WIRE_37,
		 S => SYNTHESIZED_WIRE_23,
		 C_out => SYNTHESIZED_WIRE_2);


SYNTHESIZED_WIRE_27 <= NOT(SYNTHESIZED_WIRE_35);




b2v_inst9 : full_adder
PORT MAP(A => SYNTHESIZED_WIRE_39,
		 B => SYNTHESIZED_WIRE_31,
		 C_in => SYNTHESIZED_WIRE_32,
		 S => SYNTHESIZED_WIRE_41,
		 C_out => SYNTHESIZED_WIRE_9);


END bdf_type;