-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Thu Oct 30 15:55:44 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Parte_F IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        sda : IN STD_LOGIC := '0';
        ack : OUT STD_LOGIC;
        hab_dir : OUT STD_LOGIC;
        hab_dato : OUT STD_LOGIC
    );
END Parte_F;

ARCHITECTURE BEHAVIOR OF Parte_F IS
    TYPE type_fstate IS (Guardar_dir,R_W,ACK1,Guardar_dato,Oscioso);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,fin_dir,soy,fin_dato,sda)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Oscioso;
            ack <= '0';
            hab_dir <= '0';
            hab_dato <= '0';
        ELSE
            ack <= '0';
            hab_dir <= '0';
            hab_dato <= '0';
            CASE fstate IS
                WHEN Guardar_dir =>
                    IF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= R_W;
                    ELSIF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guardar_dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardar_dir;
                    END IF;

                    hab_dato <= '0';

                    hab_dir <= '1';

                    ack <= '0';
                WHEN R_W =>
                    reg_fstate <= ACK1;

                    hab_dato <= '0';

                    hab_dir <= '0';

                    ack <= '0';
                WHEN ACK1 =>
                    reg_fstate <= Guardar_dato;

                    hab_dato <= '0';

                    hab_dir <= '0';

                    ack <= '1';
                WHEN Guardar_dato =>
                    IF ((fin_dato = '0')) THEN
                        reg_fstate <= Guardar_dato;
                    ELSIF ((fin_dato = '1')) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardar_dato;
                    END IF;

                    hab_dato <= '1';

                    hab_dir <= '0';

                    ack <= '0';
                WHEN Oscioso =>
                    IF ((sda = '1')) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((sda = '0')) THEN
                        reg_fstate <= Guardar_dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oscioso;
                    END IF;

                    hab_dato <= '0';

                    hab_dir <= '0';

                    ack <= '0';
                WHEN OTHERS => 
                    ack <= 'X';
                    hab_dir <= 'X';
                    hab_dato <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
